lab3.vhdl
